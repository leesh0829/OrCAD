** Profile: "SCHEMATIC1-ronaldo"  [ D:\Or CAD\2022 pspice dinon\rlc-PSpiceFiles\SCHEMATIC1\ronaldo.sim ] 

** Creating circuit file "ronaldo.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
* From [PSPICE NETLIST] section of C:\SPB_Data\cdssetup\OrCAD_PSpice\17.2.0\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 39ms 0 
.STEP LIN PARAM cv 0.5uF 1.5uF 0.1uF 
.OPTIONS ADVCONV
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC1.net" 


.END
